netcdf Input1 {
dimensions:
    time = 3 ;
    ID = 2 ;
variables:
    double time(time) ;
        time:units = "days since 2000-01-01 00:00:00" ;
        time:calendar = "standard" ;
    float precipitation(ID, time) ;
    int ID(ID) ;

data:
    time = 0, 1, 2 ;
    ID = 2, 1 ;
    precipitation =
         1.0, 1.1, 1.2,
         2.0, 2.1, 2.2 ;
}
