netcdf Input2 {
dimensions:
    time = 3 ;
    ID = 3 ;
variables:
    double time(time) ;
        time:units = "days since 2000-01-01 00:00:00" ;
        time:calendar = "standard" ;
    float precipitation(ID, time) ;
    int ID(ID) ;

data:
    time = 0, 1, 2 ;
    ID = 3, 4, 5 ;
    precipitation =
         3.0, 3.1, 3.2,
         4.0, 4.1, 4.2,
         5.0, 5.1, 5.2 ;
}
